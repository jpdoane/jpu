//uart

`include "jpu_defines.vh"

`define UART_PARITY 1
`define UART_DATA_WIDTH 8
`define UART_STOP_BITS 1
`define UART_DEFAULT_BAUDRATE  9600
`define UART_CLK_FREQ `CLK_FREQ  

`define UART_DIVIDE_OVERRIDE_SIM 8


