////
`define DEBUG_ON (* mark_debug = "true" *) (* KEEP = "TRUE" *) (* DONT_TOUCH = "TRUE" *)
`define DEBUG_OFF  

`define UART_DEBUG `DEBUG_OFF
`define TOP_DEBUG `DEBUG_ON
`define CORE_DEBUG `DEBUG_OFF

